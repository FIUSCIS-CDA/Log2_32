// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition"
// CREATED		"Sun Apr 27 16:27:16 2025"

module Log2_32(
	A,
	log2
);


input wire	[31:0] A;
output wire	[4:0] log2;

wire	SYNTHESIZED_WIRE_0;
wire	SYNTHESIZED_WIRE_1;
wire	SYNTHESIZED_WIRE_2;
wire	SYNTHESIZED_WIRE_3;
wire	SYNTHESIZED_WIRE_4;
wire	SYNTHESIZED_WIRE_5;
wire	SYNTHESIZED_WIRE_6;
wire	SYNTHESIZED_WIRE_7;
wire	SYNTHESIZED_WIRE_8;
wire	SYNTHESIZED_WIRE_9;
wire	SYNTHESIZED_WIRE_10;
wire	SYNTHESIZED_WIRE_11;
wire	SYNTHESIZED_WIRE_12;
wire	SYNTHESIZED_WIRE_13;
wire	SYNTHESIZED_WIRE_14;
wire	SYNTHESIZED_WIRE_15;
wire	SYNTHESIZED_WIRE_16;
wire	SYNTHESIZED_WIRE_17;
wire	SYNTHESIZED_WIRE_18;
wire	SYNTHESIZED_WIRE_19;
wire	SYNTHESIZED_WIRE_20;
wire	SYNTHESIZED_WIRE_21;
wire	SYNTHESIZED_WIRE_22;
wire	SYNTHESIZED_WIRE_23;
wire	SYNTHESIZED_WIRE_24;
wire	SYNTHESIZED_WIRE_25;
wire	SYNTHESIZED_WIRE_26;
wire	SYNTHESIZED_WIRE_27;
wire	SYNTHESIZED_WIRE_28;
wire	SYNTHESIZED_WIRE_29;
wire	SYNTHESIZED_WIRE_30;
wire	SYNTHESIZED_WIRE_122;
wire	SYNTHESIZED_WIRE_32;
wire	SYNTHESIZED_WIRE_123;
wire	SYNTHESIZED_WIRE_34;
wire	SYNTHESIZED_WIRE_124;
wire	SYNTHESIZED_WIRE_36;
wire	SYNTHESIZED_WIRE_125;
wire	SYNTHESIZED_WIRE_38;
wire	SYNTHESIZED_WIRE_126;
wire	SYNTHESIZED_WIRE_40;
wire	SYNTHESIZED_WIRE_127;
wire	SYNTHESIZED_WIRE_42;
wire	SYNTHESIZED_WIRE_128;
wire	SYNTHESIZED_WIRE_44;
wire	SYNTHESIZED_WIRE_129;
wire	SYNTHESIZED_WIRE_46;
wire	SYNTHESIZED_WIRE_130;
wire	SYNTHESIZED_WIRE_48;
wire	SYNTHESIZED_WIRE_131;
wire	SYNTHESIZED_WIRE_50;
wire	SYNTHESIZED_WIRE_132;
wire	SYNTHESIZED_WIRE_52;
wire	SYNTHESIZED_WIRE_133;
wire	SYNTHESIZED_WIRE_54;
wire	SYNTHESIZED_WIRE_134;
wire	SYNTHESIZED_WIRE_56;
wire	SYNTHESIZED_WIRE_135;
wire	SYNTHESIZED_WIRE_58;
wire	SYNTHESIZED_WIRE_136;
wire	SYNTHESIZED_WIRE_60;
wire	SYNTHESIZED_WIRE_137;
wire	SYNTHESIZED_WIRE_62;
wire	SYNTHESIZED_WIRE_138;
wire	SYNTHESIZED_WIRE_64;
wire	SYNTHESIZED_WIRE_139;
wire	SYNTHESIZED_WIRE_66;
wire	SYNTHESIZED_WIRE_140;
wire	SYNTHESIZED_WIRE_68;
wire	SYNTHESIZED_WIRE_141;
wire	SYNTHESIZED_WIRE_70;
wire	SYNTHESIZED_WIRE_142;
wire	SYNTHESIZED_WIRE_72;
wire	SYNTHESIZED_WIRE_143;
wire	SYNTHESIZED_WIRE_74;
wire	SYNTHESIZED_WIRE_144;
wire	SYNTHESIZED_WIRE_76;
wire	SYNTHESIZED_WIRE_145;
wire	SYNTHESIZED_WIRE_78;
wire	SYNTHESIZED_WIRE_146;
wire	SYNTHESIZED_WIRE_80;
wire	SYNTHESIZED_WIRE_147;
wire	SYNTHESIZED_WIRE_82;
wire	SYNTHESIZED_WIRE_148;
wire	SYNTHESIZED_WIRE_84;
wire	SYNTHESIZED_WIRE_149;
wire	SYNTHESIZED_WIRE_86;
wire	SYNTHESIZED_WIRE_150;
wire	SYNTHESIZED_WIRE_88;
wire	SYNTHESIZED_WIRE_151;
wire	SYNTHESIZED_WIRE_90;
wire	SYNTHESIZED_WIRE_121;




assign	SYNTHESIZED_WIRE_122 =  ~A[31];


Encoder_32	b2v_inst1(
	.A0(SYNTHESIZED_WIRE_0),
	.A1(SYNTHESIZED_WIRE_1),
	.A2(SYNTHESIZED_WIRE_2),
	.A3(SYNTHESIZED_WIRE_3),
	.A4(SYNTHESIZED_WIRE_4),
	.A5(SYNTHESIZED_WIRE_5),
	.A6(SYNTHESIZED_WIRE_6),
	.A7(SYNTHESIZED_WIRE_7),
	.A8(SYNTHESIZED_WIRE_8),
	.A9(SYNTHESIZED_WIRE_9),
	.A10(SYNTHESIZED_WIRE_10),
	.A11(SYNTHESIZED_WIRE_11),
	.A12(SYNTHESIZED_WIRE_12),
	.A13(SYNTHESIZED_WIRE_13),
	.A14(SYNTHESIZED_WIRE_14),
	.A15(SYNTHESIZED_WIRE_15),
	.A16(SYNTHESIZED_WIRE_16),
	.A17(SYNTHESIZED_WIRE_17),
	.A18(SYNTHESIZED_WIRE_18),
	.A19(SYNTHESIZED_WIRE_19),
	.A20(SYNTHESIZED_WIRE_20),
	.A21(SYNTHESIZED_WIRE_21),
	.A22(SYNTHESIZED_WIRE_22),
	.A23(SYNTHESIZED_WIRE_23),
	.A24(SYNTHESIZED_WIRE_24),
	.A25(SYNTHESIZED_WIRE_25),
	.A26(SYNTHESIZED_WIRE_26),
	.A27(SYNTHESIZED_WIRE_27),
	.A28(SYNTHESIZED_WIRE_28),
	.A29(SYNTHESIZED_WIRE_29),
	.A30(SYNTHESIZED_WIRE_30),
	.A31(A[31]),
	.Q(log2));

assign	SYNTHESIZED_WIRE_48 =  ~A[22];

assign	SYNTHESIZED_WIRE_50 =  ~A[21];

assign	SYNTHESIZED_WIRE_123 = SYNTHESIZED_WIRE_122 & SYNTHESIZED_WIRE_32;

assign	SYNTHESIZED_WIRE_52 =  ~A[20];

assign	SYNTHESIZED_WIRE_54 =  ~A[19];

assign	SYNTHESIZED_WIRE_56 =  ~A[18];

assign	SYNTHESIZED_WIRE_58 =  ~A[17];

assign	SYNTHESIZED_WIRE_60 =  ~A[16];

assign	SYNTHESIZED_WIRE_62 =  ~A[15];

assign	SYNTHESIZED_WIRE_32 =  ~A[30];

assign	SYNTHESIZED_WIRE_64 =  ~A[14];

assign	SYNTHESIZED_WIRE_66 =  ~A[13];

assign	SYNTHESIZED_WIRE_124 = SYNTHESIZED_WIRE_123 & SYNTHESIZED_WIRE_34;

assign	SYNTHESIZED_WIRE_125 = SYNTHESIZED_WIRE_124 & SYNTHESIZED_WIRE_36;

assign	SYNTHESIZED_WIRE_68 =  ~A[12];

assign	SYNTHESIZED_WIRE_70 =  ~A[11];

assign	SYNTHESIZED_WIRE_72 =  ~A[10];

assign	SYNTHESIZED_WIRE_74 =  ~A[9];

assign	SYNTHESIZED_WIRE_76 =  ~A[8];

assign	SYNTHESIZED_WIRE_78 =  ~A[7];

assign	SYNTHESIZED_WIRE_34 =  ~A[29];

assign	SYNTHESIZED_WIRE_80 =  ~A[6];

assign	SYNTHESIZED_WIRE_82 =  ~A[5];

assign	SYNTHESIZED_WIRE_84 =  ~A[4];

assign	SYNTHESIZED_WIRE_86 =  ~A[3];

assign	SYNTHESIZED_WIRE_88 =  ~A[2];

assign	SYNTHESIZED_WIRE_90 =  ~A[1];

assign	SYNTHESIZED_WIRE_126 = SYNTHESIZED_WIRE_125 & SYNTHESIZED_WIRE_38;

assign	SYNTHESIZED_WIRE_127 = SYNTHESIZED_WIRE_126 & SYNTHESIZED_WIRE_40;

assign	SYNTHESIZED_WIRE_128 = SYNTHESIZED_WIRE_127 & SYNTHESIZED_WIRE_42;

assign	SYNTHESIZED_WIRE_129 = SYNTHESIZED_WIRE_128 & SYNTHESIZED_WIRE_44;

assign	SYNTHESIZED_WIRE_36 =  ~A[28];

assign	SYNTHESIZED_WIRE_130 = SYNTHESIZED_WIRE_129 & SYNTHESIZED_WIRE_46;

assign	SYNTHESIZED_WIRE_131 = SYNTHESIZED_WIRE_130 & SYNTHESIZED_WIRE_48;

assign	SYNTHESIZED_WIRE_132 = SYNTHESIZED_WIRE_131 & SYNTHESIZED_WIRE_50;

assign	SYNTHESIZED_WIRE_133 = SYNTHESIZED_WIRE_132 & SYNTHESIZED_WIRE_52;

assign	SYNTHESIZED_WIRE_134 = SYNTHESIZED_WIRE_133 & SYNTHESIZED_WIRE_54;

assign	SYNTHESIZED_WIRE_135 = SYNTHESIZED_WIRE_134 & SYNTHESIZED_WIRE_56;

assign	SYNTHESIZED_WIRE_136 = SYNTHESIZED_WIRE_135 & SYNTHESIZED_WIRE_58;

assign	SYNTHESIZED_WIRE_137 = SYNTHESIZED_WIRE_136 & SYNTHESIZED_WIRE_60;

assign	SYNTHESIZED_WIRE_138 = SYNTHESIZED_WIRE_137 & SYNTHESIZED_WIRE_62;

assign	SYNTHESIZED_WIRE_139 = SYNTHESIZED_WIRE_138 & SYNTHESIZED_WIRE_64;

assign	SYNTHESIZED_WIRE_38 =  ~A[27];

assign	SYNTHESIZED_WIRE_140 = SYNTHESIZED_WIRE_139 & SYNTHESIZED_WIRE_66;

assign	SYNTHESIZED_WIRE_141 = SYNTHESIZED_WIRE_140 & SYNTHESIZED_WIRE_68;

assign	SYNTHESIZED_WIRE_142 = SYNTHESIZED_WIRE_141 & SYNTHESIZED_WIRE_70;

assign	SYNTHESIZED_WIRE_143 = SYNTHESIZED_WIRE_142 & SYNTHESIZED_WIRE_72;

assign	SYNTHESIZED_WIRE_144 = SYNTHESIZED_WIRE_143 & SYNTHESIZED_WIRE_74;

assign	SYNTHESIZED_WIRE_145 = SYNTHESIZED_WIRE_144 & SYNTHESIZED_WIRE_76;

assign	SYNTHESIZED_WIRE_146 = SYNTHESIZED_WIRE_145 & SYNTHESIZED_WIRE_78;

assign	SYNTHESIZED_WIRE_147 = SYNTHESIZED_WIRE_146 & SYNTHESIZED_WIRE_80;

assign	SYNTHESIZED_WIRE_148 = SYNTHESIZED_WIRE_147 & SYNTHESIZED_WIRE_82;

assign	SYNTHESIZED_WIRE_149 = SYNTHESIZED_WIRE_148 & SYNTHESIZED_WIRE_84;

assign	SYNTHESIZED_WIRE_40 =  ~A[26];

assign	SYNTHESIZED_WIRE_150 = SYNTHESIZED_WIRE_149 & SYNTHESIZED_WIRE_86;

assign	SYNTHESIZED_WIRE_151 = SYNTHESIZED_WIRE_150 & SYNTHESIZED_WIRE_88;

assign	SYNTHESIZED_WIRE_121 = SYNTHESIZED_WIRE_151 & SYNTHESIZED_WIRE_90;

assign	SYNTHESIZED_WIRE_30 = SYNTHESIZED_WIRE_122 & A[30];

assign	SYNTHESIZED_WIRE_29 = SYNTHESIZED_WIRE_123 & A[29];

assign	SYNTHESIZED_WIRE_28 = SYNTHESIZED_WIRE_124 & A[28];

assign	SYNTHESIZED_WIRE_27 = SYNTHESIZED_WIRE_125 & A[27];

assign	SYNTHESIZED_WIRE_26 = SYNTHESIZED_WIRE_126 & A[26];

assign	SYNTHESIZED_WIRE_25 = SYNTHESIZED_WIRE_127 & A[25];

assign	SYNTHESIZED_WIRE_24 = SYNTHESIZED_WIRE_128 & A[24];

assign	SYNTHESIZED_WIRE_42 =  ~A[25];

assign	SYNTHESIZED_WIRE_23 = SYNTHESIZED_WIRE_129 & A[23];

assign	SYNTHESIZED_WIRE_22 = SYNTHESIZED_WIRE_130 & A[22];

assign	SYNTHESIZED_WIRE_21 = SYNTHESIZED_WIRE_131 & A[21];

assign	SYNTHESIZED_WIRE_20 = SYNTHESIZED_WIRE_132 & A[20];

assign	SYNTHESIZED_WIRE_19 = SYNTHESIZED_WIRE_133 & A[19];

assign	SYNTHESIZED_WIRE_18 = SYNTHESIZED_WIRE_134 & A[18];

assign	SYNTHESIZED_WIRE_17 = SYNTHESIZED_WIRE_135 & A[17];

assign	SYNTHESIZED_WIRE_16 = SYNTHESIZED_WIRE_136 & A[16];

assign	SYNTHESIZED_WIRE_15 = SYNTHESIZED_WIRE_137 & A[15];

assign	SYNTHESIZED_WIRE_14 = SYNTHESIZED_WIRE_138 & A[14];

assign	SYNTHESIZED_WIRE_44 =  ~A[24];

assign	SYNTHESIZED_WIRE_13 = SYNTHESIZED_WIRE_139 & A[13];

assign	SYNTHESIZED_WIRE_12 = SYNTHESIZED_WIRE_140 & A[12];

assign	SYNTHESIZED_WIRE_11 = SYNTHESIZED_WIRE_141 & A[11];

assign	SYNTHESIZED_WIRE_10 = SYNTHESIZED_WIRE_142 & A[10];

assign	SYNTHESIZED_WIRE_9 = SYNTHESIZED_WIRE_143 & A[9];

assign	SYNTHESIZED_WIRE_8 = SYNTHESIZED_WIRE_144 & A[8];

assign	SYNTHESIZED_WIRE_7 = SYNTHESIZED_WIRE_145 & A[7];

assign	SYNTHESIZED_WIRE_6 = SYNTHESIZED_WIRE_146 & A[6];

assign	SYNTHESIZED_WIRE_5 = SYNTHESIZED_WIRE_147 & A[5];

assign	SYNTHESIZED_WIRE_4 = SYNTHESIZED_WIRE_148 & A[4];

assign	SYNTHESIZED_WIRE_46 =  ~A[23];

assign	SYNTHESIZED_WIRE_3 = SYNTHESIZED_WIRE_149 & A[3];

assign	SYNTHESIZED_WIRE_2 = SYNTHESIZED_WIRE_150 & A[2];

assign	SYNTHESIZED_WIRE_1 = SYNTHESIZED_WIRE_151 & A[1];

assign	SYNTHESIZED_WIRE_0 = SYNTHESIZED_WIRE_121 & A[0];


endmodule
